version https://git-lfs.github.com/spec/v1
oid sha256:3e894a667773208b7e063f3fcd5fb343c2bbdc752dd00bdc450534138ac9af81
size 19341
