version https://git-lfs.github.com/spec/v1
oid sha256:31918258c405cb9c54c1ca8eb86c172a1fd94c9a346f83635fc9e7d2792b10c5
size 359349
