version https://git-lfs.github.com/spec/v1
oid sha256:bb5ca91725a2fcf0bc723e4d4dc3ee8292486486db80c2fbaf5104c6401581df
size 10258
