version https://git-lfs.github.com/spec/v1
oid sha256:8bb96003a1175e604fbce9a54e9a012a323aaab969cfb2d61bd054788a7906eb
size 9641
