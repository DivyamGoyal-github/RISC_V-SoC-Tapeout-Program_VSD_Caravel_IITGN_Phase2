version https://git-lfs.github.com/spec/v1
oid sha256:2f0e79878049b2f0121ac038d401d51b5191e6bed5299ddc6f2631a10ec2f1d4
size 98735678
